library ieee;
use ieee.std_logic_1164.all;

entity light_flasher is
--  Port ( );
end light_flasher;

architecture behavioral_light_flasher of light_flasher is

begin


end behavioral_light_flasher;
