library ieee;
use ieee.std_logic_1164.all;

entity bootstrapper is
    -- TODO: implement
end;

architecture behavioral_bootstrapper of bootstrapper is
    -- TODO: implement
begin
end;
